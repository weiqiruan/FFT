module cf_fft_1024_8_6 (clock_c, i1, i2, i3, i4, i5, o1, o2, o3);
input  clock_c;
input  i1;
input  [15:0] i2;
input  [15:0] i3;
input  i4;
input  i5;
output o1;
output [15:0] o2;
output [15:0] o3;
wire   s1_1;
wire   [15:0] s1_2;
wire   [15:0] s1_3;
wire   s2_1;
wire   [15:0] s2_2;
wire   [15:0] s2_3;
wire   s3_1;
wire   [15:0] s3_2;
wire   [15:0] s3_3;
wire   s4_1;
wire   [15:0] s4_2;
wire   [15:0] s4_3;
wire   s5_1;
wire   [15:0] s5_2;
wire   [15:0] s5_3;
wire   s6_1;
wire   [15:0] s6_2;
wire   [15:0] s6_3;
wire   s7_1;
wire   [15:0] s7_2;
wire   [15:0] s7_3;
wire   s8_1;
wire   [15:0] s8_2;
wire   [15:0] s8_3;
cf_fft_1024_8_21 s1 (clock_c, s2_1, s2_2, s2_3, i4, i5, s1_1, s1_2, s1_3);
cf_fft_1024_8_19 s2 (clock_c, s3_1, s3_2, s3_3, i4, i5, s2_1, s2_2, s2_3);
cf_fft_1024_8_17 s3 (clock_c, s4_1, s4_2, s4_3, i4, i5, s3_1, s3_2, s3_3);
cf_fft_1024_8_15 s4 (clock_c, s5_1, s5_2, s5_3, i4, i5, s4_1, s4_2, s4_3);
cf_fft_1024_8_13 s5 (clock_c, s6_1, s6_2, s6_3, i4, i5, s5_1, s5_2, s5_3);
cf_fft_1024_8_11 s6 (clock_c, s7_1, s7_2, s7_3, i4, i5, s6_1, s6_2, s6_3);
cf_fft_1024_8_9 s7 (clock_c, s8_1, s8_2, s8_3, i4, i5, s7_1, s7_2, s7_3);
cf_fft_1024_8_7 s8 (clock_c, i1, i2, i3, i4, i5, s8_1, s8_2, s8_3);
assign o3 = s1_3;
assign o2 = s1_2;
assign o1 = s1_1;
endmodule
