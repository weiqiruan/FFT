module cf_fft_1024_8 (clock_c, enable_i, reset_i, sync_i, data_0_i, data_1_i, sync_o, data_0_o, data_1_o);
input  clock_c;
input  enable_i;
input  reset_i;
input  sync_i;
input  [15:0] data_0_i;
input  [15:0] data_1_i;
output sync_o;
output [15:0] data_0_o;
output [15:0] data_1_o;
wire   n1;
wire   [15:0] n2;
wire   [15:0] n3;
cf_fft_1024_8_1 s1 (clock_c, sync_i, data_0_i, data_1_i, enable_i, reset_i, n1, n2, n3);
assign sync_o = n1;
assign data_0_o = n2;
assign data_1_o = n3;
endmodule

module cf_fft_1024_8_1 (clock_c, i1, i2, i3, i4, i5, o1, o2, o3);
input  clock_c;
input  i1;
input  [15:0] i2;
input  [15:0] i3;
input  i4;
input  i5;
output o1;
output [15:0] o2;
output [15:0] o3;
wire   s1_1;
wire   [15:0] s1_2;
wire   [15:0] s1_3;
wire   s2_1;
wire   [15:0] s2_2;
wire   [15:0] s2_3;
wire   s3_1;
wire   [15:0] s3_2;
wire   [15:0] s3_3;
wire   s4_1;
wire   [15:0] s4_2;
wire   [15:0] s4_3;
cf_fft_1024_8_23 s1 (clock_c, s3_1, s3_2, s3_3, i4, i5, s1_1, s1_2, s1_3);
cf_fft_1024_8_6 s2 (clock_c, s1_1, s1_2, s1_3, i4, i5, s2_1, s2_2, s2_3);
cf_fft_1024_8_5 s3 (clock_c, s4_1, s4_2, s4_3, i4, i5, s3_1, s3_2, s3_3);
cf_fft_1024_8_2 s4 (clock_c, i1, i2, i3, i4, i5, s4_1, s4_2, s4_3);
assign o3 = s2_3;
assign o2 = s2_2;
assign o1 = s2_1;
endmodule
