module cf_fft_1024_8_37 (i1, i2, i3, i4, i5, i6, i7, i8, o1);
input  i1;
input  i2;
input  i3;
input  i4;
input  i5;
input  i6;
input  i7;
input  [2:0] i8;
output o1;
wire   [2:0] n1;
wire   [2:0] n2;
wire   [2:0] n3;
wire   n4;
wire   n5;
wire   n6;
wire   n7;
wire   n8;
wire   n9;
wire   s10_1;
assign n1 = 3'b010;
assign n2 = 3'b100;
assign n3 = 3'b110;
assign n4 = i8 == n1;
assign n5 = i8 == n2;
assign n6 = i8 == n3;
assign n7 = n6 ? i5 : s10_1;
assign n8 = n5 ? i6 : n7;
assign n9 = n4 ? i7 : n8;
cf_fft_1024_8_38 s10 (i1, i2, i3, i4, i8, s10_1);
assign o1 = n9;
endmodule
