module cf_fft_1024_8_22 (clock_c, i1, i2, i3, i4, i5, o1, o2);
input  clock_c;
input  [15:0] i1;
input  [15:0] i2;
input  [8:0] i3;
input  i4;
input  i5;
output [15:0] o1;
output [15:0] o2;
reg    [15:0] n1;
wire   [7:0] n2;
wire   [7:0] n3;
reg    [15:0] n4;
wire   [7:0] n5;
wire   [7:0] n6;
reg    [7:0] n7;
reg    [7:0] n8;
reg    [7:0] n9;
reg    [7:0] n10;
reg    [15:0] n11;
wire   [7:0] n12;
wire   [7:0] n13;
wire   [15:0] n14;
wire   [7:0] n15;
reg    [7:0] n16;
wire   [15:0] n17;
wire   [7:0] n18;
reg    [7:0] n19;
wire   [7:0] n20;
reg    [7:0] n21;
wire   [15:0] n22;
wire   [7:0] n23;
reg    [7:0] n24;
wire   [15:0] n25;
wire   [7:0] n26;
reg    [7:0] n27;
wire   [7:0] n28;
reg    [7:0] n29;
wire   [7:0] n30;
wire   [7:0] n31;
wire   [15:0] n32;
reg    [15:0] n33;
wire   [7:0] n34;
wire   [7:0] n35;
wire   [15:0] n36;
reg    [15:0] n37;
initial n1 = 16'b0000000000000000;
always @ (posedge clock_c)
  if (i5 == 1'b1)
    n1 <= 16'b0000000000000000;
  else if (i4 == 1'b1)
    n1 <= i1;
assign n2 = {n1[15],
  n1[14],
  n1[13],
  n1[12],
  n1[11],
  n1[10],
  n1[9],
  n1[8]};
assign n3 = {n1[7],
  n1[6],
  n1[5],
  n1[4],
  n1[3],
  n1[2],
  n1[1],
  n1[0]};
initial n4 = 16'b0000000000000000;
always @ (posedge clock_c)
  if (i5 == 1'b1)
    n4 <= 16'b0000000000000000;
  else if (i4 == 1'b1)
    n4 <= i2;
assign n5 = {n4[15],
  n4[14],
  n4[13],
  n4[12],
  n4[11],
  n4[10],
  n4[9],
  n4[8]};
assign n6 = {n4[7],
  n4[6],
  n4[5],
  n4[4],
  n4[3],
  n4[2],
  n4[1],
  n4[0]};
initial n7 = 8'b00000000;
always @ (posedge clock_c)
  if (i5 == 1'b1)
    n7 <= 8'b00000000;
  else if (i4 == 1'b1)
    n7 <= n2;
initial n8 = 8'b00000000;
always @ (posedge clock_c)
  if (i5 == 1'b1)
    n8 <= 8'b00000000;
  else if (i4 == 1'b1)
    n8 <= n7;
initial n9 = 8'b00000000;
always @ (posedge clock_c)
  if (i5 == 1'b1)
    n9 <= 8'b00000000;
  else if (i4 == 1'b1)
    n9 <= n3;
initial n10 = 8'b00000000;
always @ (posedge clock_c)
  if (i5 == 1'b1)
    n10 <= 8'b00000000;
  else if (i4 == 1'b1)
    n10 <= n9;
initial n11 = 16'b0000000000000000;
always @ (posedge clock_c)
  if (i4 == 1'b1)
    case (i3)
      9'b000000000 : n11 <= 16'b0111111100000000;
      9'b000000001 : n11 <= 16'b0111111111111111;
      9'b000000010 : n11 <= 16'b0111111111111110;
      9'b000000011 : n11 <= 16'b0111111111111101;
      9'b000000100 : n11 <= 16'b0111111111111100;
      9'b000000101 : n11 <= 16'b0111111111111100;
      9'b000000110 : n11 <= 16'b0111111111111011;
      9'b000000111 : n11 <= 16'b0111111111111010;
      9'b000001000 : n11 <= 16'b0111111111111001;
      9'b000001001 : n11 <= 16'b0111111111111000;
      9'b000001010 : n11 <= 16'b0111111111111000;
      9'b000001011 : n11 <= 16'b0111111111110111;
      9'b000001100 : n11 <= 16'b0111111111110110;
      9'b000001101 : n11 <= 16'b0111111111110101;
      9'b000001110 : n11 <= 16'b0111111111110101;
      9'b000001111 : n11 <= 16'b0111111111110100;
      9'b000010000 : n11 <= 16'b0111111111110011;
      9'b000010001 : n11 <= 16'b0111111111110010;
      9'b000010010 : n11 <= 16'b0111111111110001;
      9'b000010011 : n11 <= 16'b0111111111110001;
      9'b000010100 : n11 <= 16'b0111111111110000;
      9'b000010101 : n11 <= 16'b0111111011101111;
      9'b000010110 : n11 <= 16'b0111111011101110;
      9'b000010111 : n11 <= 16'b0111111011101101;
      9'b000011000 : n11 <= 16'b0111111011101101;
      9'b000011001 : n11 <= 16'b0111111011101100;
      9'b000011010 : n11 <= 16'b0111111011101011;
      9'b000011011 : n11 <= 16'b0111111011101010;
      9'b000011100 : n11 <= 16'b0111111011101010;
      9'b000011101 : n11 <= 16'b0111110111101001;
      9'b000011110 : n11 <= 16'b0111110111101000;
      9'b000011111 : n11 <= 16'b0111110111100111;
      9'b000100000 : n11 <= 16'b0111110111100111;
      9'b000100001 : n11 <= 16'b0111110111100110;
      9'b000100010 : n11 <= 16'b0111110111100101;
      9'b000100011 : n11 <= 16'b0111110111100100;
      9'b000100100 : n11 <= 16'b0111110011100011;
      9'b000100101 : n11 <= 16'b0111110011100011;
      9'b000100110 : n11 <= 16'b0111110011100010;
      9'b000100111 : n11 <= 16'b0111110011100001;
      9'b000101000 : n11 <= 16'b0111110011100000;
      9'b000101001 : n11 <= 16'b0111101111100000;
      9'b000101010 : n11 <= 16'b0111101111011111;
      9'b000101011 : n11 <= 16'b0111101111011110;
      9'b000101100 : n11 <= 16'b0111101111011101;
      9'b000101101 : n11 <= 16'b0111101111011101;
      9'b000101110 : n11 <= 16'b0111101011011100;
      9'b000101111 : n11 <= 16'b0111101011011011;
      9'b000110000 : n11 <= 16'b0111101011011010;
      9'b000110001 : n11 <= 16'b0111101011011010;
      9'b000110010 : n11 <= 16'b0111101011011001;
      9'b000110011 : n11 <= 16'b0111100111011000;
      9'b000110100 : n11 <= 16'b0111100111010111;
      9'b000110101 : n11 <= 16'b0111100111010111;
      9'b000110110 : n11 <= 16'b0111100111010110;
      9'b000110111 : n11 <= 16'b0111100011010101;
      9'b000111000 : n11 <= 16'b0111100011010100;
      9'b000111001 : n11 <= 16'b0111100011010100;
      9'b000111010 : n11 <= 16'b0111011111010011;
      9'b000111011 : n11 <= 16'b0111011111010010;
      9'b000111100 : n11 <= 16'b0111011111010001;
      9'b000111101 : n11 <= 16'b0111011111010001;
      9'b000111110 : n11 <= 16'b0111011011010000;
      9'b000111111 : n11 <= 16'b0111011011001111;
      9'b001000000 : n11 <= 16'b0111011011001111;
      9'b001000001 : n11 <= 16'b0111010111001110;
      9'b001000010 : n11 <= 16'b0111010111001101;
      9'b001000011 : n11 <= 16'b0111010111001100;
      9'b001000100 : n11 <= 16'b0111010111001100;
      9'b001000101 : n11 <= 16'b0111010011001011;
      9'b001000110 : n11 <= 16'b0111010011001010;
      9'b001000111 : n11 <= 16'b0111010011001001;
      9'b001001000 : n11 <= 16'b0111001111001001;
      9'b001001001 : n11 <= 16'b0111001111001000;
      9'b001001010 : n11 <= 16'b0111001111000111;
      9'b001001011 : n11 <= 16'b0111001011000111;
      9'b001001100 : n11 <= 16'b0111001011000110;
      9'b001001101 : n11 <= 16'b0111000111000101;
      9'b001001110 : n11 <= 16'b0111000111000101;
      9'b001001111 : n11 <= 16'b0111000111000100;
      9'b001010000 : n11 <= 16'b0111000011000011;
      9'b001010001 : n11 <= 16'b0111000011000010;
      9'b001010010 : n11 <= 16'b0111000011000010;
      9'b001010011 : n11 <= 16'b0110111111000001;
      9'b001010100 : n11 <= 16'b0110111111000000;
      9'b001010101 : n11 <= 16'b0110111011000000;
      9'b001010110 : n11 <= 16'b0110111010111111;
      9'b001010111 : n11 <= 16'b0110111010111110;
      9'b001011000 : n11 <= 16'b0110110110111110;
      9'b001011001 : n11 <= 16'b0110110110111101;
      9'b001011010 : n11 <= 16'b0110110010111100;
      9'b001011011 : n11 <= 16'b0110110010111100;
      9'b001011100 : n11 <= 16'b0110110010111011;
      9'b001011101 : n11 <= 16'b0110101110111010;
      9'b001011110 : n11 <= 16'b0110101110111010;
      9'b001011111 : n11 <= 16'b0110101010111001;
      9'b001100000 : n11 <= 16'b0110101010111000;
      9'b001100001 : n11 <= 16'b0110100110111000;
      9'b001100010 : n11 <= 16'b0110100110110111;
      9'b001100011 : n11 <= 16'b0110100110110110;
      9'b001100100 : n11 <= 16'b0110100010110110;
      9'b001100101 : n11 <= 16'b0110100010110101;
      9'b001100110 : n11 <= 16'b0110011110110101;
      9'b001100111 : n11 <= 16'b0110011110110100;
      9'b001101000 : n11 <= 16'b0110011010110011;
      9'b001101001 : n11 <= 16'b0110011010110011;
      9'b001101010 : n11 <= 16'b0110010110110010;
      9'b001101011 : n11 <= 16'b0110010110110001;
      9'b001101100 : n11 <= 16'b0110010010110001;
      9'b001101101 : n11 <= 16'b0110010010110000;
      9'b001101110 : n11 <= 16'b0110001110110000;
      9'b001101111 : n11 <= 16'b0110001110101111;
      9'b001110000 : n11 <= 16'b0110001010101110;
      9'b001110001 : n11 <= 16'b0110001010101110;
      9'b001110010 : n11 <= 16'b0110000110101101;
      9'b001110011 : n11 <= 16'b0110000110101100;
      9'b001110100 : n11 <= 16'b0110000010101100;
      9'b001110101 : n11 <= 16'b0110000010101011;
      9'b001110110 : n11 <= 16'b0101111110101011;
      9'b001110111 : n11 <= 16'b0101111110101010;
      9'b001111000 : n11 <= 16'b0101111010101010;
      9'b001111001 : n11 <= 16'b0101111010101001;
      9'b001111010 : n11 <= 16'b0101110110101000;
      9'b001111011 : n11 <= 16'b0101110110101000;
      9'b001111100 : n11 <= 16'b0101110010100111;
      9'b001111101 : n11 <= 16'b0101110010100111;
      9'b001111110 : n11 <= 16'b0101101110100110;
      9'b001111111 : n11 <= 16'b0101101110100110;
      9'b010000000 : n11 <= 16'b0101101010100101;
      9'b010000001 : n11 <= 16'b0101100110100100;
      9'b010000010 : n11 <= 16'b0101100110100100;
      9'b010000011 : n11 <= 16'b0101100010100011;
      9'b010000100 : n11 <= 16'b0101100010100011;
      9'b010000101 : n11 <= 16'b0101011110100010;
      9'b010000110 : n11 <= 16'b0101011110100010;
      9'b010000111 : n11 <= 16'b0101011010100001;
      9'b010001000 : n11 <= 16'b0101010110100001;
      9'b010001001 : n11 <= 16'b0101010110100000;
      9'b010001010 : n11 <= 16'b0101010010100000;
      9'b010001011 : n11 <= 16'b0101010010011111;
      9'b010001100 : n11 <= 16'b0101001110011111;
      9'b010001101 : n11 <= 16'b0101001110011110;
      9'b010001110 : n11 <= 16'b0101001010011110;
      9'b010001111 : n11 <= 16'b0101000110011101;
      9'b010010000 : n11 <= 16'b0101000110011101;
      9'b010010001 : n11 <= 16'b0101000010011100;
      9'b010010010 : n11 <= 16'b0100111110011100;
      9'b010010011 : n11 <= 16'b0100111110011011;
      9'b010010100 : n11 <= 16'b0100111010011011;
      9'b010010101 : n11 <= 16'b0100111010011010;
      9'b010010110 : n11 <= 16'b0100110110011010;
      9'b010010111 : n11 <= 16'b0100110010011001;
      9'b010011000 : n11 <= 16'b0100110010011001;
      9'b010011001 : n11 <= 16'b0100101110011000;
      9'b010011010 : n11 <= 16'b0100101010011000;
      9'b010011011 : n11 <= 16'b0100101010010111;
      9'b010011100 : n11 <= 16'b0100100110010111;
      9'b010011101 : n11 <= 16'b0100100110010110;
      9'b010011110 : n11 <= 16'b0100100010010110;
      9'b010011111 : n11 <= 16'b0100011110010110;
      9'b010100000 : n11 <= 16'b0100011110010101;
      9'b010100001 : n11 <= 16'b0100011010010101;
      9'b010100010 : n11 <= 16'b0100010110010100;
      9'b010100011 : n11 <= 16'b0100010110010100;
      9'b010100100 : n11 <= 16'b0100010010010011;
      9'b010100101 : n11 <= 16'b0100001110010011;
      9'b010100110 : n11 <= 16'b0100001110010011;
      9'b010100111 : n11 <= 16'b0100001010010010;
      9'b010101000 : n11 <= 16'b0100000110010010;
      9'b010101001 : n11 <= 16'b0100000110010001;
      9'b010101010 : n11 <= 16'b0100000010010001;
      9'b010101011 : n11 <= 16'b0011111110010001;
      9'b010101100 : n11 <= 16'b0011111110010000;
      9'b010101101 : n11 <= 16'b0011111010010000;
      9'b010101110 : n11 <= 16'b0011110110001111;
      9'b010101111 : n11 <= 16'b0011110110001111;
      9'b010110000 : n11 <= 16'b0011110010001111;
      9'b010110001 : n11 <= 16'b0011101110001110;
      9'b010110010 : n11 <= 16'b0011101010001110;
      9'b010110011 : n11 <= 16'b0011101010001110;
      9'b010110100 : n11 <= 16'b0011100110001101;
      9'b010110101 : n11 <= 16'b0011100010001101;
      9'b010110110 : n11 <= 16'b0011100010001100;
      9'b010110111 : n11 <= 16'b0011011110001100;
      9'b010111000 : n11 <= 16'b0011011010001100;
      9'b010111001 : n11 <= 16'b0011011010001011;
      9'b010111010 : n11 <= 16'b0011010110001011;
      9'b010111011 : n11 <= 16'b0011010010001011;
      9'b010111100 : n11 <= 16'b0011001110001010;
      9'b010111101 : n11 <= 16'b0011001110001010;
      9'b010111110 : n11 <= 16'b0011001010001010;
      9'b010111111 : n11 <= 16'b0011000110001010;
      9'b011000000 : n11 <= 16'b0011000010001001;
      9'b011000001 : n11 <= 16'b0011000010001001;
      9'b011000010 : n11 <= 16'b0010111110001001;
      9'b011000011 : n11 <= 16'b0010111010001000;
      9'b011000100 : n11 <= 16'b0010111010001000;
      9'b011000101 : n11 <= 16'b0010110110001000;
      9'b011000110 : n11 <= 16'b0010110010001000;
      9'b011000111 : n11 <= 16'b0010101110000111;
      9'b011001000 : n11 <= 16'b0010101110000111;
      9'b011001001 : n11 <= 16'b0010101010000111;
      9'b011001010 : n11 <= 16'b0010100110000110;
      9'b011001011 : n11 <= 16'b0010100010000110;
      9'b011001100 : n11 <= 16'b0010100010000110;
      9'b011001101 : n11 <= 16'b0010011110000110;
      9'b011001110 : n11 <= 16'b0010011010000101;
      9'b011001111 : n11 <= 16'b0010010110000101;
      9'b011010000 : n11 <= 16'b0010010110000101;
      9'b011010001 : n11 <= 16'b0010010010000101;
      9'b011010010 : n11 <= 16'b0010001110000101;
      9'b011010011 : n11 <= 16'b0010001010000100;
      9'b011010100 : n11 <= 16'b0010001010000100;
      9'b011010101 : n11 <= 16'b0010000110000100;
      9'b011010110 : n11 <= 16'b0010000010000100;
      9'b011010111 : n11 <= 16'b0001111110000100;
      9'b011011000 : n11 <= 16'b0001111110000011;
      9'b011011001 : n11 <= 16'b0001111010000011;
      9'b011011010 : n11 <= 16'b0001110110000011;
      9'b011011011 : n11 <= 16'b0001110010000011;
      9'b011011100 : n11 <= 16'b0001110010000011;
      9'b011011101 : n11 <= 16'b0001101110000010;
      9'b011011110 : n11 <= 16'b0001101010000010;
      9'b011011111 : n11 <= 16'b0001100110000010;
      9'b011100000 : n11 <= 16'b0001100010000010;
      9'b011100001 : n11 <= 16'b0001100010000010;
      9'b011100010 : n11 <= 16'b0001011110000010;
      9'b011100011 : n11 <= 16'b0001011010000010;
      9'b011100100 : n11 <= 16'b0001010110000001;
      9'b011100101 : n11 <= 16'b0001010110000001;
      9'b011100110 : n11 <= 16'b0001010010000001;
      9'b011100111 : n11 <= 16'b0001001110000001;
      9'b011101000 : n11 <= 16'b0001001010000001;
      9'b011101001 : n11 <= 16'b0001001010000001;
      9'b011101010 : n11 <= 16'b0001000110000001;
      9'b011101011 : n11 <= 16'b0001000010000001;
      9'b011101100 : n11 <= 16'b0000111110000000;
      9'b011101101 : n11 <= 16'b0000111010000000;
      9'b011101110 : n11 <= 16'b0000111010000000;
      9'b011101111 : n11 <= 16'b0000110110000000;
      9'b011110000 : n11 <= 16'b0000110010000000;
      9'b011110001 : n11 <= 16'b0000101110000000;
      9'b011110010 : n11 <= 16'b0000101010000000;
      9'b011110011 : n11 <= 16'b0000101010000000;
      9'b011110100 : n11 <= 16'b0000100110000000;
      9'b011110101 : n11 <= 16'b0000100010000000;
      9'b011110110 : n11 <= 16'b0000011110000000;
      9'b011110111 : n11 <= 16'b0000011110000000;
      9'b011111000 : n11 <= 16'b0000011010000000;
      9'b011111001 : n11 <= 16'b0000010110000000;
      9'b011111010 : n11 <= 16'b0000010010000000;
      9'b011111011 : n11 <= 16'b0000001110000000;
      9'b011111100 : n11 <= 16'b0000001110000000;
      9'b011111101 : n11 <= 16'b0000001010000000;
      9'b011111110 : n11 <= 16'b0000000110000000;
      9'b011111111 : n11 <= 16'b0000000010000000;
      9'b100000000 : n11 <= 16'b0000000010000000;
      9'b100000001 : n11 <= 16'b1111111110000000;
      9'b100000010 : n11 <= 16'b1111111010000000;
      9'b100000011 : n11 <= 16'b1111110110000000;
      9'b100000100 : n11 <= 16'b1111110010000000;
      9'b100000101 : n11 <= 16'b1111110010000000;
      9'b100000110 : n11 <= 16'b1111101110000000;
      9'b100000111 : n11 <= 16'b1111101010000000;
      9'b100001000 : n11 <= 16'b1111100110000000;
      9'b100001001 : n11 <= 16'b1111100010000000;
      9'b100001010 : n11 <= 16'b1111100010000000;
      9'b100001011 : n11 <= 16'b1111011110000000;
      9'b100001100 : n11 <= 16'b1111011010000000;
      9'b100001101 : n11 <= 16'b1111010110000000;
      9'b100001110 : n11 <= 16'b1111010110000000;
      9'b100001111 : n11 <= 16'b1111010010000000;
      9'b100010000 : n11 <= 16'b1111001110000000;
      9'b100010001 : n11 <= 16'b1111001010000000;
      9'b100010010 : n11 <= 16'b1111000110000000;
      9'b100010011 : n11 <= 16'b1111000110000000;
      9'b100010100 : n11 <= 16'b1111000010000000;
      9'b100010101 : n11 <= 16'b1110111110000001;
      9'b100010110 : n11 <= 16'b1110111010000001;
      9'b100010111 : n11 <= 16'b1110110110000001;
      9'b100011000 : n11 <= 16'b1110110110000001;
      9'b100011001 : n11 <= 16'b1110110010000001;
      9'b100011010 : n11 <= 16'b1110101110000001;
      9'b100011011 : n11 <= 16'b1110101010000001;
      9'b100011100 : n11 <= 16'b1110101010000001;
      9'b100011101 : n11 <= 16'b1110100110000010;
      9'b100011110 : n11 <= 16'b1110100010000010;
      9'b100011111 : n11 <= 16'b1110011110000010;
      9'b100100000 : n11 <= 16'b1110011110000010;
      9'b100100001 : n11 <= 16'b1110011010000010;
      9'b100100010 : n11 <= 16'b1110010110000010;
      9'b100100011 : n11 <= 16'b1110010010000010;
      9'b100100100 : n11 <= 16'b1110001110000011;
      9'b100100101 : n11 <= 16'b1110001110000011;
      9'b100100110 : n11 <= 16'b1110001010000011;
      9'b100100111 : n11 <= 16'b1110000110000011;
      9'b100101000 : n11 <= 16'b1110000010000011;
      9'b100101001 : n11 <= 16'b1110000010000100;
      9'b100101010 : n11 <= 16'b1101111110000100;
      9'b100101011 : n11 <= 16'b1101111010000100;
      9'b100101100 : n11 <= 16'b1101110110000100;
      9'b100101101 : n11 <= 16'b1101110110000100;
      9'b100101110 : n11 <= 16'b1101110010000101;
      9'b100101111 : n11 <= 16'b1101101110000101;
      9'b100110000 : n11 <= 16'b1101101010000101;
      9'b100110001 : n11 <= 16'b1101101010000101;
      9'b100110010 : n11 <= 16'b1101100110000101;
      9'b100110011 : n11 <= 16'b1101100010000110;
      9'b100110100 : n11 <= 16'b1101011110000110;
      9'b100110101 : n11 <= 16'b1101011110000110;
      9'b100110110 : n11 <= 16'b1101011010000110;
      9'b100110111 : n11 <= 16'b1101010110000111;
      9'b100111000 : n11 <= 16'b1101010010000111;
      9'b100111001 : n11 <= 16'b1101010010000111;
      9'b100111010 : n11 <= 16'b1101001110001000;
      9'b100111011 : n11 <= 16'b1101001010001000;
      9'b100111100 : n11 <= 16'b1101000110001000;
      9'b100111101 : n11 <= 16'b1101000110001000;
      9'b100111110 : n11 <= 16'b1101000010001001;
      9'b100111111 : n11 <= 16'b1100111110001001;
      9'b101000000 : n11 <= 16'b1100111110001001;
      9'b101000001 : n11 <= 16'b1100111010001010;
      9'b101000010 : n11 <= 16'b1100110110001010;
      9'b101000011 : n11 <= 16'b1100110010001010;
      9'b101000100 : n11 <= 16'b1100110010001010;
      9'b101000101 : n11 <= 16'b1100101110001011;
      9'b101000110 : n11 <= 16'b1100101010001011;
      9'b101000111 : n11 <= 16'b1100100110001011;
      9'b101001000 : n11 <= 16'b1100100110001100;
      9'b101001001 : n11 <= 16'b1100100010001100;
      9'b101001010 : n11 <= 16'b1100011110001100;
      9'b101001011 : n11 <= 16'b1100011110001101;
      9'b101001100 : n11 <= 16'b1100011010001101;
      9'b101001101 : n11 <= 16'b1100010110001110;
      9'b101001110 : n11 <= 16'b1100010110001110;
      9'b101001111 : n11 <= 16'b1100010010001110;
      9'b101010000 : n11 <= 16'b1100001110001111;
      9'b101010001 : n11 <= 16'b1100001010001111;
      9'b101010010 : n11 <= 16'b1100001010001111;
      9'b101010011 : n11 <= 16'b1100000110010000;
      9'b101010100 : n11 <= 16'b1100000010010000;
      9'b101010101 : n11 <= 16'b1100000010010001;
      9'b101010110 : n11 <= 16'b1011111110010001;
      9'b101010111 : n11 <= 16'b1011111010010001;
      9'b101011000 : n11 <= 16'b1011111010010010;
      9'b101011001 : n11 <= 16'b1011110110010010;
      9'b101011010 : n11 <= 16'b1011110010010011;
      9'b101011011 : n11 <= 16'b1011110010010011;
      9'b101011100 : n11 <= 16'b1011101110010011;
      9'b101011101 : n11 <= 16'b1011101010010100;
      9'b101011110 : n11 <= 16'b1011101010010100;
      9'b101011111 : n11 <= 16'b1011100110010101;
      9'b101100000 : n11 <= 16'b1011100010010101;
      9'b101100001 : n11 <= 16'b1011100010010110;
      9'b101100010 : n11 <= 16'b1011011110010110;
      9'b101100011 : n11 <= 16'b1011011010010110;
      9'b101100100 : n11 <= 16'b1011011010010111;
      9'b101100101 : n11 <= 16'b1011010110010111;
      9'b101100110 : n11 <= 16'b1011010110011000;
      9'b101100111 : n11 <= 16'b1011010010011000;
      9'b101101000 : n11 <= 16'b1011001110011001;
      9'b101101001 : n11 <= 16'b1011001110011001;
      9'b101101010 : n11 <= 16'b1011001010011010;
      9'b101101011 : n11 <= 16'b1011000110011010;
      9'b101101100 : n11 <= 16'b1011000110011011;
      9'b101101101 : n11 <= 16'b1011000010011011;
      9'b101101110 : n11 <= 16'b1011000010011100;
      9'b101101111 : n11 <= 16'b1010111110011100;
      9'b101110000 : n11 <= 16'b1010111010011101;
      9'b101110001 : n11 <= 16'b1010111010011101;
      9'b101110010 : n11 <= 16'b1010110110011110;
      9'b101110011 : n11 <= 16'b1010110010011110;
      9'b101110100 : n11 <= 16'b1010110010011111;
      9'b101110101 : n11 <= 16'b1010101110011111;
      9'b101110110 : n11 <= 16'b1010101110100000;
      9'b101110111 : n11 <= 16'b1010101010100000;
      9'b101111000 : n11 <= 16'b1010101010100001;
      9'b101111001 : n11 <= 16'b1010100110100001;
      9'b101111010 : n11 <= 16'b1010100010100010;
      9'b101111011 : n11 <= 16'b1010100010100010;
      9'b101111100 : n11 <= 16'b1010011110100011;
      9'b101111101 : n11 <= 16'b1010011110100011;
      9'b101111110 : n11 <= 16'b1010011010100100;
      9'b101111111 : n11 <= 16'b1010011010100100;
      9'b110000000 : n11 <= 16'b1010010110100101;
      9'b110000001 : n11 <= 16'b1010010010100110;
      9'b110000010 : n11 <= 16'b1010010010100110;
      9'b110000011 : n11 <= 16'b1010001110100111;
      9'b110000100 : n11 <= 16'b1010001110100111;
      9'b110000101 : n11 <= 16'b1010001010101000;
      9'b110000110 : n11 <= 16'b1010001010101000;
      9'b110000111 : n11 <= 16'b1010000110101001;
      9'b110001000 : n11 <= 16'b1010000110101010;
      9'b110001001 : n11 <= 16'b1010000010101010;
      9'b110001010 : n11 <= 16'b1010000010101011;
      9'b110001011 : n11 <= 16'b1001111110101011;
      9'b110001100 : n11 <= 16'b1001111110101100;
      9'b110001101 : n11 <= 16'b1001111010101100;
      9'b110001110 : n11 <= 16'b1001111010101101;
      9'b110001111 : n11 <= 16'b1001110110101110;
      9'b110010000 : n11 <= 16'b1001110110101110;
      9'b110010001 : n11 <= 16'b1001110010101111;
      9'b110010010 : n11 <= 16'b1001110010110000;
      9'b110010011 : n11 <= 16'b1001101110110000;
      9'b110010100 : n11 <= 16'b1001101110110001;
      9'b110010101 : n11 <= 16'b1001101010110001;
      9'b110010110 : n11 <= 16'b1001101010110010;
      9'b110010111 : n11 <= 16'b1001100110110011;
      9'b110011000 : n11 <= 16'b1001100110110011;
      9'b110011001 : n11 <= 16'b1001100010110100;
      9'b110011010 : n11 <= 16'b1001100010110101;
      9'b110011011 : n11 <= 16'b1001011110110101;
      9'b110011100 : n11 <= 16'b1001011110110110;
      9'b110011101 : n11 <= 16'b1001011010110110;
      9'b110011110 : n11 <= 16'b1001011010110111;
      9'b110011111 : n11 <= 16'b1001011010111000;
      9'b110100000 : n11 <= 16'b1001010110111000;
      9'b110100001 : n11 <= 16'b1001010110111001;
      9'b110100010 : n11 <= 16'b1001010010111010;
      9'b110100011 : n11 <= 16'b1001010010111010;
      9'b110100100 : n11 <= 16'b1001001110111011;
      9'b110100101 : n11 <= 16'b1001001110111100;
      9'b110100110 : n11 <= 16'b1001001110111100;
      9'b110100111 : n11 <= 16'b1001001010111101;
      9'b110101000 : n11 <= 16'b1001001010111110;
      9'b110101001 : n11 <= 16'b1001000110111110;
      9'b110101010 : n11 <= 16'b1001000110111111;
      9'b110101011 : n11 <= 16'b1001000111000000;
      9'b110101100 : n11 <= 16'b1001000011000000;
      9'b110101101 : n11 <= 16'b1001000011000001;
      9'b110101110 : n11 <= 16'b1000111111000010;
      9'b110101111 : n11 <= 16'b1000111111000010;
      9'b110110000 : n11 <= 16'b1000111111000011;
      9'b110110001 : n11 <= 16'b1000111011000100;
      9'b110110010 : n11 <= 16'b1000111011000101;
      9'b110110011 : n11 <= 16'b1000111011000101;
      9'b110110100 : n11 <= 16'b1000110111000110;
      9'b110110101 : n11 <= 16'b1000110111000111;
      9'b110110110 : n11 <= 16'b1000110011000111;
      9'b110110111 : n11 <= 16'b1000110011001000;
      9'b110111000 : n11 <= 16'b1000110011001001;
      9'b110111001 : n11 <= 16'b1000101111001001;
      9'b110111010 : n11 <= 16'b1000101111001010;
      9'b110111011 : n11 <= 16'b1000101111001011;
      9'b110111100 : n11 <= 16'b1000101011001100;
      9'b110111101 : n11 <= 16'b1000101011001100;
      9'b110111110 : n11 <= 16'b1000101011001101;
      9'b110111111 : n11 <= 16'b1000101011001110;
      9'b111000000 : n11 <= 16'b1000100111001111;
      9'b111000001 : n11 <= 16'b1000100111001111;
      9'b111000010 : n11 <= 16'b1000100111010000;
      9'b111000011 : n11 <= 16'b1000100011010001;
      9'b111000100 : n11 <= 16'b1000100011010001;
      9'b111000101 : n11 <= 16'b1000100011010010;
      9'b111000110 : n11 <= 16'b1000100011010011;
      9'b111000111 : n11 <= 16'b1000011111010100;
      9'b111001000 : n11 <= 16'b1000011111010100;
      9'b111001001 : n11 <= 16'b1000011111010101;
      9'b111001010 : n11 <= 16'b1000011011010110;
      9'b111001011 : n11 <= 16'b1000011011010111;
      9'b111001100 : n11 <= 16'b1000011011010111;
      9'b111001101 : n11 <= 16'b1000011011011000;
      9'b111001110 : n11 <= 16'b1000010111011001;
      9'b111001111 : n11 <= 16'b1000010111011010;
      9'b111010000 : n11 <= 16'b1000010111011010;
      9'b111010001 : n11 <= 16'b1000010111011011;
      9'b111010010 : n11 <= 16'b1000010111011100;
      9'b111010011 : n11 <= 16'b1000010011011101;
      9'b111010100 : n11 <= 16'b1000010011011101;
      9'b111010101 : n11 <= 16'b1000010011011110;
      9'b111010110 : n11 <= 16'b1000010011011111;
      9'b111010111 : n11 <= 16'b1000010011100000;
      9'b111011000 : n11 <= 16'b1000001111100000;
      9'b111011001 : n11 <= 16'b1000001111100001;
      9'b111011010 : n11 <= 16'b1000001111100010;
      9'b111011011 : n11 <= 16'b1000001111100011;
      9'b111011100 : n11 <= 16'b1000001111100011;
      9'b111011101 : n11 <= 16'b1000001011100100;
      9'b111011110 : n11 <= 16'b1000001011100101;
      9'b111011111 : n11 <= 16'b1000001011100110;
      9'b111100000 : n11 <= 16'b1000001011100111;
      9'b111100001 : n11 <= 16'b1000001011100111;
      9'b111100010 : n11 <= 16'b1000001011101000;
      9'b111100011 : n11 <= 16'b1000001011101001;
      9'b111100100 : n11 <= 16'b1000000111101010;
      9'b111100101 : n11 <= 16'b1000000111101010;
      9'b111100110 : n11 <= 16'b1000000111101011;
      9'b111100111 : n11 <= 16'b1000000111101100;
      9'b111101000 : n11 <= 16'b1000000111101101;
      9'b111101001 : n11 <= 16'b1000000111101101;
      9'b111101010 : n11 <= 16'b1000000111101110;
      9'b111101011 : n11 <= 16'b1000000111101111;
      9'b111101100 : n11 <= 16'b1000000011110000;
      9'b111101101 : n11 <= 16'b1000000011110001;
      9'b111101110 : n11 <= 16'b1000000011110001;
      9'b111101111 : n11 <= 16'b1000000011110010;
      9'b111110000 : n11 <= 16'b1000000011110011;
      9'b111110001 : n11 <= 16'b1000000011110100;
      9'b111110010 : n11 <= 16'b1000000011110101;
      9'b111110011 : n11 <= 16'b1000000011110101;
      9'b111110100 : n11 <= 16'b1000000011110110;
      9'b111110101 : n11 <= 16'b1000000011110111;
      9'b111110110 : n11 <= 16'b1000000011111000;
      9'b111110111 : n11 <= 16'b1000000011111000;
      9'b111111000 : n11 <= 16'b1000000011111001;
      9'b111111001 : n11 <= 16'b1000000011111010;
      9'b111111010 : n11 <= 16'b1000000011111011;
      9'b111111011 : n11 <= 16'b1000000011111100;
      9'b111111100 : n11 <= 16'b1000000011111100;
      9'b111111101 : n11 <= 16'b1000000011111101;
      9'b111111110 : n11 <= 16'b1000000011111110;
      9'b111111111 : n11 <= 16'b1000000011111111;
      default : n11 <= 16'bxxxxxxxxxxxxxxxx;
    endcase
assign n12 = {n11[15],
  n11[14],
  n11[13],
  n11[12],
  n11[11],
  n11[10],
  n11[9],
  n11[8]};
assign n13 = {n11[7],
  n11[6],
  n11[5],
  n11[4],
  n11[3],
  n11[2],
  n11[1],
  n11[0]};
assign n14 = {{8{n5[7]}}, n5} * {{8{n12[7]}}, n12};
assign n15 = {n14[14],
  n14[13],
  n14[12],
  n14[11],
  n14[10],
  n14[9],
  n14[8],
  n14[7]};
initial n16 = 8'b00000000;
always @ (posedge clock_c)
  if (i5 == 1'b1)
    n16 <= 8'b00000000;
  else if (i4 == 1'b1)
    n16 <= n15;
assign n17 = {{8{n6[7]}}, n6} * {{8{n13[7]}}, n13};
assign n18 = {n17[14],
  n17[13],
  n17[12],
  n17[11],
  n17[10],
  n17[9],
  n17[8],
  n17[7]};
initial n19 = 8'b00000000;
always @ (posedge clock_c)
  if (i5 == 1'b1)
    n19 <= 8'b00000000;
  else if (i4 == 1'b1)
    n19 <= n18;
assign n20 = n16 - n19;
initial n21 = 8'b00000000;
always @ (posedge clock_c)
  if (i5 == 1'b1)
    n21 <= 8'b00000000;
  else if (i4 == 1'b1)
    n21 <= n20;
assign n22 = {{8{n5[7]}}, n5} * {{8{n13[7]}}, n13};
assign n23 = {n22[14],
  n22[13],
  n22[12],
  n22[11],
  n22[10],
  n22[9],
  n22[8],
  n22[7]};
initial n24 = 8'b00000000;
always @ (posedge clock_c)
  if (i5 == 1'b1)
    n24 <= 8'b00000000;
  else if (i4 == 1'b1)
    n24 <= n23;
assign n25 = {{8{n6[7]}}, n6} * {{8{n12[7]}}, n12};
assign n26 = {n25[14],
  n25[13],
  n25[12],
  n25[11],
  n25[10],
  n25[9],
  n25[8],
  n25[7]};
initial n27 = 8'b00000000;
always @ (posedge clock_c)
  if (i5 == 1'b1)
    n27 <= 8'b00000000;
  else if (i4 == 1'b1)
    n27 <= n26;
assign n28 = n24 + n27;
initial n29 = 8'b00000000;
always @ (posedge clock_c)
  if (i5 == 1'b1)
    n29 <= 8'b00000000;
  else if (i4 == 1'b1)
    n29 <= n28;
assign n30 = n8 + n21;
assign n31 = n10 + n29;
assign n32 = {n30, n31};
initial n33 = 16'b0000000000000000;
always @ (posedge clock_c)
  if (i5 == 1'b1)
    n33 <= 16'b0000000000000000;
  else if (i4 == 1'b1)
    n33 <= n32;
assign n34 = n8 - n21;
assign n35 = n10 - n29;
assign n36 = {n34, n35};
initial n37 = 16'b0000000000000000;
always @ (posedge clock_c)
  if (i5 == 1'b1)
    n37 <= 16'b0000000000000000;
  else if (i4 == 1'b1)
    n37 <= n36;
assign o2 = n37;
assign o1 = n33;
endmodule
