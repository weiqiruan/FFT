module cf_fft_1024_8_36 (o1, o2, o3, o4, o5, o6, o7, o8);
output o1;
output o2;
output o3;
output o4;
output o5;
output o6;
output o7;
output o8;
wire   n1;
wire   n2;
wire   n3;
wire   n4;
wire   n5;
wire   n6;
wire   n7;
wire   n8;
assign n1 = 1'b0;
assign n2 = 1'b1;
assign n3 = 1'b0;
assign n4 = 1'b1;
assign n5 = 1'b0;
assign n6 = 1'b1;
assign n7 = 1'b0;
assign n8 = 1'b0;
assign o8 = n8;
assign o7 = n7;
assign o6 = n6;
assign o5 = n5;
assign o4 = n4;
assign o3 = n3;
assign o2 = n2;
assign o1 = n1;
endmodule
